
package metro_mpi_pkg;

parameter CREDIT_WIDTH = 3;

//typedef logic [63:0]  reg64_t;


/*typedef enum logic [1:0] {
    ENUM1  = 2'b00,
    ENUM2  = 2'b01,
    ENUM3  = 2'b10,
    ENUM3  = 2'b11
} enum_name;    // Enum*/



endpackage
